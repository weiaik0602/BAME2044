library verilog;
use verilog.vl_types.all;
entity Integrate_tb is
end Integrate_tb;

library verilog;
use verilog.vl_types.all;
entity lab_dp_tb is
    generic(
        S0              : integer := 0;
        S1              : integer := 1;
        S2              : integer := 2;
        S3              : integer := 8;
        S4              : integer := 9;
        S5              : integer := 10;
        S6              : integer := 11;
        S7              : integer := 12;
        S8              : integer := 13;
        S9              : integer := 14;
        S10             : integer := 15
    );
end lab_dp_tb;
